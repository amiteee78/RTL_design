`timescale 1ns/1ns
`include "apb_arch.svh"

module apb_mem (apbif.mem membus);

endmodule